module pipeline_unit (
    input  wire         clk,
    input  wire         reset,
    input  wire [31:0]  inputs,
    input  wire         in_valid,
    input  wire         flush,
    output wire [31:0]  outputs, 
    output wire         out_valid
);

// actual pipeline stages here

// stage 1

// stage 2

// stage ...


endmodule