`include "defines.vh"

module consumer (
    input  wire clk,
    input  wire reset,

    input  wire [`DATA_WIDTH-1:0] in_data,
    input  wire [`ID_WIDTH-1:0]   in_id,
    input  wire                   in_valid
);
// Consumer logic placeholder
endmodule