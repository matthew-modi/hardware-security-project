module buffer_slots (
    input  wire        clk,
    input  wire        reset,
    input  wire [31:0] inputs,
    input  wire        stall,
    output wire [31:0] outputs,
    output wire        to_stall_mgmt
);
    // Stall and Regular Slots 
endmodule
