module arbiter (
    input  wire clk,
    input  wire reset,
    input  wire req_1,
    input  wire req_2,
    output wire grant_1,
    output wire grant_2
);
// Arbitration logic placeholder
endmodule