`define PIPELINE_DEPTH 3

`define ADDRESS_WIDTH 8
`define DATA_WIDTH 32
`define ID_WIDTH 8

`define RESOURCE_DELAY 10
`define RESOURCE_DELAY_COUNTER_WIDTH 4