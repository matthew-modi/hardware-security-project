module arbiter (
    input  wire clk,
    input  wire reset,

    input  wire in_valid_1,
    input  wire in_valid_2,

    output wire out_stall_1,
    output wire out_stall_2
);
// Arbitration logic placeholder
endmodule